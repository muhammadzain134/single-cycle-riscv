`timescale 1ns / 1ps

module ALU_control(
input logic [6:0] funct7,
input logic [2:0] finct3,
input logic [1:0] ALUOp,
output logic [3:0] control_sig
    );
    
    always_comb begin
        case(ALUOp)
            2'b00: 
                control_sig = 4'b0000;
            2'b01:
                control_sig = 4'b1000;
            2'b10:  // R-type
                case(finct3)
                3'b000: 
                    if(funct7[5]== 0)
                        control_sig = 4'b0000; // Add
                    else
                        control_sig = 4'b1000; // Sub
                3'b001: control_sig = 4'b0001; // shift left logical
                3'b010: control_sig = 4'b0010; // set less than
                3'b011: control_sig = 4'b0011; // set less than unsigned
                3'b100: control_sig = 4'b0100; // xor
                3'b101: 
                    if(funct7[5]==0)
                        control_sig = 4'b0101; // Shift right logical
                    else
                        control_sig = 4'b1101; // Shift right arithmatic
                3'b110: control_sig = 4'b0110; // or
                3'b111: control_sig = 4'b0111; // and
                endcase
            2'b11: // I-type
                case(finct3)
                3'b000: control_sig = 4'b0000;
                3'b001: control_sig = 4'b0001;
                3'b010: control_sig = 4'b0010;
                3'b011: control_sig = 4'b0011;
                3'b100: control_sig = 4'b0100;
                3'b101: 
                    if(funct7[5]==0)
                        control_sig = 4'b0101; // Shift right logical immediate
                    else
                        control_sig = 4'b1101; // Shift right arithmatic immediate
                3'b110: control_sig = 4'b0110;
                3'b111: control_sig = 4'b0111;
                 endcase
              default:  control_sig = 4'b1111; 
        endcase
    
    end

endmodule
